// $Id: $
// File name:   tb_ATD_block.sv
// Created:     12/4/2017
// Author:      Kartikeya Mishra
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: test bench for the overall atd block



`timescale 1ns/100 ps

module tb_ATD_block();
	
	localparam NUM_CNT_BITS = 8;
	localparam CLK_PERIOD = 2.5;

	reg tb_clk;
	//reg tb_atd_clock;
	reg tb_n_rst;
	reg tb_ATD_data;
	reg tb_ATD_clk;
	
	reg tb_data_taken;
	reg tb_data_ready;
	reg [127:0] tb_ATD_parallel;
	
	
	
	// Clock generation block
	always
	begin
		tb_clk = 1'b0;
		#(CLK_PERIOD/2.0);
		tb_clk = 1'b1;
		#(CLK_PERIOD/2.0);
	end

	//DUT map port
	ATD_block DUT(.clk(tb_clk), .n_rst(tb_n_rst), .ATD_data(tb_ATD_data), .ATD_clk(tb_ATD_clk), .data_taken(tb_data_taken), .data_ready(tb_data_ready), .ATD_parallel(tb_ATD_parallel));

	initial begin
		tb_n_rst = 1'b0;
		tb_ATD_data = 1'b1;
		tb_ATD_clk = 1'b0;
		
		tb_data_taken = '0;
		
		@(posedge tb_clk);
		@(posedge tb_clk);

		//test case 1: checking for data 
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_ATD_data = '0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		tb_ATD_data = '1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		tb_ATD_data = '0;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_ATD_data = '1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_ATD_data = '0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_ATD_data = '1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		tb_ATD_data = '0;
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;		
		@(posedge tb_clk); 
		@(posedge tb_clk);
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	

		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;		
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		

		tb_ATD_clk = 1'b1;			
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	

		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	

		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		@(posedge tb_clk); 
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		tb_n_rst 	= 1'b1;
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);
		tb_ATD_clk = 1'b1;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b0;
		@(posedge tb_clk);
		@(posedge tb_clk);		
		tb_ATD_clk = 1'b1;	
		if(tb_data_ready == '1)  begin
			$info("data_ready working !!");
		end
		else
		begin
			$error("data ready not working");
		end
end

/*task task_name;
	input  input;
begin
	//Task stuff
end
endtask*/
endmodule	
